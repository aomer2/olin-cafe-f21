module shift_left_logical(in, shamt, out);

parameter N = 32; // only used as a constant! Don't feel like you need to a shifter for arbitrary N.

input wire [N-1:0] in;            // the input number that will be shifted left. Fill in the remainder with zeros.
input wire [$clog2(N)-1:0] shamt; // the amount to shift by (think of it as a decimal number from 0 to 31). 
output logic [N-1:0] out; 

always_comb begin : left_shift
    out = 0;

    for (int i = 0; i < N; i = i + 1) begin
        if ((i + shamt) < N) out[i + shamt] = in[i];
    end

end


endmodule
